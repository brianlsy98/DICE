* delay_line with switch_cap_inverters

.subckt delay_line_combination_1 gnd vdd vin vout
* first stage inv
MP0  vin_bar  vin      vdd   vdd  pmos  W='MP0W'  L='MP0L'
MN0  vin_bar  vin      gnd   gnd  nmos  W='MN0W'  L='MN0L'
MN4  vin_bar  VCTRL_1  mn4s  gnd  nmos  W='MN4W'  L='MN4L'
C0   mn4s     gnd      'C0'
C1   vin_bar  gnd      'C1'
* second stage inv
MP1  vin_bb   vin_bar  vdd   vdd  pmos  W='MP1W'  L='MP1L'
MN1  vin_bb   vin_bar  gnd   gnd  nmos  W='MN1W'  L='MN1L'
MN5  vin_bb   VCTRL_2  mn5s  gnd  nmos  W='MN5W'  L='MN5L'
C2   mn5s     gnd      'C2'
C3   vin_bb   gnd      'C3'
* third stage inv
MP2  vout_b   vin_bb   vdd   vdd  pmos  W='MP2W'  L='MP2L'
MN2  vout_b   vin_bb   gnd   gnd  nmos  W='MN2W'  L='MN2L'
MN6  vout_b   VCTRL_2  mn6s  gnd  nmos  W='MN6W'  L='MN6L'
C4   mn6s     gnd      'C4'
C5   vout_b   gnd      'C5'
* fourth stage inv
MP3  vout     vout_b   vdd   vdd  pmos  W='MP3W'  L='MP3L'
MN3  vout     vout_b   gnd   gnd  nmos  W='MN3W'  L='MN3L'
C7   vout     gnd      'C7'
* vctrls
VCTRL_1 VCTRL_1 0 'VCTRL_1'
VCTRL_2 VCTRL_2 0 'VCTRL_2'
VCTRL_3 VCTRL_3 0 'VCTRL_3'
.ends delay_line_combination_1