* Tan_CLIA_Pin_3 Amplifier

.subckt tan_clia_pin_3_amp gnd vdd vinn vinp vout

* PMOS Transistors
MP0   net5   dm_1   vdd   vdd   pmos W='MP0W'  L='MP0L'
MP1   net3   net050 vdd   vdd   pmos W='MP1W'  L='MP1L'
MP2   dm_1   dm_1   vdd   vdd   pmos W='MP2W'  L='MP2L'
MP3   vout   net050 vdd   vdd   pmos W='MP3W'  L='MP3L'
MP4   net050 voutn  vdd   vdd   pmos W='MP4W'  L='MP4L'
MP5   voutn  voutn  vdd   vdd   pmos W='MP5W'  L='MP5L'
MP6   net8   vinp   net31 net31 pmos W='MP6W'  L='MP6L'
MP7   dm_2   vinn   net31 net31 pmos W='MP7W'  L='MP7L'
MP8   net31  net1   vdd   vdd   pmos W='MP8W'  L='MP8L'
MP9   vb3    net1   vdd   vdd   pmos W='MP9W'  L='MP9L'
MP10  vb4    net1   vdd   vdd   pmos W='MP10W' L='MP10L'
MP11  net1   net1   vdd   vdd   pmos W='MP11W' L='MP11L'

* NMOS Transistors
MN0   net5   net3 gnd  gnd nmos W='MN0W'  L='MN0L'
MN1   net3   vb4  gnd  gnd nmos W='MN1W'  L='MN1L'
MN2   net3   net3 gnd  gnd nmos W='MN2W'  L='MN2L'
MN3   dm_2   vb4  gnd  gnd nmos W='MN3W'  L='MN3L'
MN4   voutn  vb3  dm_2 gnd nmos W='MN4W'  L='MN4L'
MN5   net8   vb4  gnd  gnd nmos W='MN5W'  L='MN5L'
MN6   net050 vb3  net8 gnd nmos W='MN6W'  L='MN6L'
MN7   net7   vb4  gnd  gnd nmos W='MN7W'  L='MN7L'
MN8   vb4    vb3  net6 gnd nmos W='MN8W'  L='MN8L'
MN9   dm_1   vb3  net7 gnd nmos W='MN9W'  L='MN9L'
MN10  net6   vb4  gnd  gnd nmos W='MN10W' L='MN10L'
MN11  vout   net5 gnd  gnd nmos W='MN11W' L='MN11L'
MN12  vb3    vb3  gnd  gnd nmos W='MN12W' L='MN12L'

* Current Source
I0 net1 gnd 'I0'

* Capacitors and Resistor
C1 net8 vout 'C1'
C0 net2 gnd 'C0'
R0 net5 net2 'R0'

.ends tan_clia_pin_3_amp
