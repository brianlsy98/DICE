* Sau_CFCC_Pin_3 Amplifier

.subckt sau_cfcc_pin_3_amp gnd vdd vinn vinp vout

* PMOS Transistors
MP0   VOUT    net050 vdd vdd pmos W='MP0W'    L='MP0L'
MP1   net049  VOUTN  vdd vdd pmos W='MP1W'    L='MP1L'
MP2   net043  net050 vdd vdd pmos W='MP2W'    L='MP2L'
MP3   net050  VOUTN  vdd vdd pmos W='MP3W'    L='MP3L'
MP4   VOUTN   VOUTN  vdd vdd pmos W='MP4W'    L='MP4L'
MP5   net063  VINP   net31 net31 pmos W='MP5W'  L='MP5L'
MP6   DM_2    VINN   net31 net31 pmos W='MP6W'  L='MP6L'
MP7   net31   net013 vdd vdd pmos W='MP7W'    L='MP7L'
MP8   VB3     net013 vdd vdd pmos W='MP8W'    L='MP8L'
MP9   DM_1    net013 vdd vdd pmos W='MP9W'    L='MP9L'
MP10  VB4     net013 vdd vdd pmos W='MP10W'   L='MP10L'
MP11  net013  net013 vdd vdd pmos W='MP11W'   L='MP11L'

* NMOS Transistors
MN0   VOUT    net049 gnd gnd nmos W='MN0W'    L='MN0L'
MN1   net049  net043 gnd gnd nmos W='MN1W'    L='MN1L'
MN2   net043  net043 gnd gnd nmos W='MN2W'    L='MN2L'
MN3   DM_2    VB4    gnd gnd nmos W='MN3W'    L='MN3L'
MN4   VOUTN   VB3    DM_2 gnd nmos W='MN4W'    L='MN4L'
MN5   net063  VB4    gnd gnd nmos W='MN5W'    L='MN5L'
MN6   net050  VB3    net063 gnd nmos W='MN6W'  L='MN6L'
MN7   net54   VB4    gnd gnd nmos W='MN7W'    L='MN7L'
MN8   VB3     VB3    gnd gnd nmos W='MN8W'    L='MN8L'
MN9   VB4     VB3    net54 gnd nmos W='MN9W'  L='MN9L'
MN10  net56   VB4    gnd gnd nmos W='MN10W'   L='MN10L'
MN11  DM_1    VB3    net56 gnd nmos W='MN11W' L='MN11L'

* Current Source
I0 net013 gnd 'CURRENT_0_BIAS'

* Capacitor
C0 net063 vout 'CAPACITOR_0'

.ends sau_cfcc_pin_3_amp
