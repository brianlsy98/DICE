* Peng_TCFC_Pin_3 Amplifier

.subckt peng_tcfc_pin_3_amp gnd vdd vinn vinp vout

MP0   net10   vb2     net049 vdd pmos W='MP0W'    L='MP0L'
MP1   vout    voutp   vdd    vdd pmos W='MP1W'    L='MP1L'
MP2   net049  vb1     vdd    vdd pmos W='MP2W'    L='MP2L'
MP3   net043  voutp   vdd    vdd pmos W='MP3W'    L='MP3L'
MP4   vb1     vb2     net2   vdd pmos W='MP4W'    L='MP4L'
MP5   vb2     vb2     vdd    vdd pmos W='MP5W'    L='MP5L'
MP6   voutp   voutn   vdd    vdd pmos W='MP6W'    L='MP6L'
MP7   voutn   voutn   vdd    vdd pmos W='MP7W'    L='MP7L'
MP8   net063  vinp    net31  net31 pmos W='MP8W'  L='MP8L'
MP9   dm_2    vinn    net31  net31 pmos W='MP9W'  L='MP9L'
MP10  net31   vb1     vdd    vdd pmos W='MP10W'   L='MP10L'
MP11  vb3     vb2     net8   vdd pmos W='MP11W'   L='MP11L'
MP12  net8    vb1     vdd    vdd pmos W='MP12W'   L='MP12L'
MP13  net7    vb2     net6   vdd pmos W='MP13W'   L='MP13L'
MP14  net6    vb1     vdd    vdd pmos W='MP14W'   L='MP14L'
MP15  vb4     vb2     net3   vdd pmos W='MP15W'   L='MP15L'
MP16  net3    vb1     vdd    vdd pmos W='MP16W'   L='MP16L'
MP17  net2    vb1     vdd    vdd pmos W='MP17W'   L='MP17L'

MN0   vout    net10   gnd    gnd nmos W='MN0W'    L='MN0L'
MN1   net043  net043  gnd    gnd nmos W='MN1W'    L='MN1L'
MN2   net10   net043  gnd    gnd nmos W='MN2W'    L='MN2L'
MN3   dm_2    vb4     gnd    gnd nmos W='MN3W'    L='MN3L'
MN4   voutn   vb3     dm_2   gnd nmos W='MN4W'    L='MN4L'
MN5   net063  vb4     gnd    gnd nmos W='MN5W'    L='MN5L'
MN6   voutp   vb3     net063 gnd nmos W='MN6W'    L='MN6L'
MN7   net54   vb4     gnd    gnd nmos W='MN7W'    L='MN7L'
MN8   vb3     vb3     gnd    gnd nmos W='MN8W'    L='MN8L'
MN9   vb4     vb3     net54  gnd nmos W='MN9W'    L='MN9L'
MN10  net56   vb4     gnd    gnd nmos W='MN10W'   L='MN10L'
MN11  net7    vb3     net56  gnd nmos W='MN11W'   L='MN11L'
MN12  net9    vb4     gnd    gnd nmos W='MN12W'   L='MN12L'
MN13  vb2     vb3     net9   gnd nmos W='MN13W'   L='MN13L'

I0    vb1     gnd     'I0'
C1    net049  vout    'C1'
C0    voutp   vout    'C0'

.ends peng_tcfc_pin_3_amp
