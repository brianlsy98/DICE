* Leung_DFCFC2_Pin_3 Amplifier

.subckt leung_dfcfc2_pin_3_amp gnd vdd vinn vinp vout
MP0   VOUT    net050 vdd vdd pmos W='MP0W'    L='MP0L'
MP1   net049  net1   vdd vdd pmos W='MP1W'    L='MP1L'
MP2   net043  net050 vdd vdd pmos W='MP2W'    L='MP2L'
MP3   net2    net050 vdd vdd pmos W='MP3W'    L='MP3L'
MP4   net050  VOUTN  vdd vdd pmos W='MP4W'    L='MP4L'
MP5   VOUTN   VOUTN  vdd vdd pmos W='MP5W'    L='MP5L'
MP6   net063  VINP   net31 net31 pmos W='MP6W'    L='MP6L'
MP7   DM_2    VINN   net31 net31 pmos W='MP7W'    L='MP7L'
MP8   net31   net1   vdd vdd pmos W='MP8W'    L='MP8L'
MP9   VB3     net1   vdd vdd pmos W='MP9W'    L='MP9L'
MP10  DM_1    net1   vdd vdd pmos W='MP10W'   L='MP10L'
MP11  VB4     net1   vdd vdd pmos W='MP11W'   L='MP11L'
MP12  net1    net1   vdd vdd pmos W='MP12W'   L='MP12L'
MN0   VOUT    net049 gnd gnd nmos W='MN0W'    L='MN0L'
MN1   net049  net043 gnd gnd nmos W='MN1W'    L='MN1L'
MN2   net043  net043 gnd gnd nmos W='MN2W'    L='MN2L'
MN3   DM_2    VB4    gnd gnd nmos W='MN3W'    L='MN3L'
MN4   VOUTN   VB3    DM_2 gnd nmos W='MN4W'   L='MN4L'
MN5   net063  VB4    gnd gnd nmos W='MN5W'    L='MN5L'
MN6   net050  VB3    net063 gnd nmos W='MN6W'   L='MN6L'
MN7   net54   VB4    gnd gnd nmos W='MN7W'    L='MN7L'
MN8   net2    VB4    gnd gnd nmos W='MN8W'    L='MN8L'
MN9   VB3     VB3    gnd gnd nmos W='MN9W'    L='MN9L'
MN10  VB4     VB3    net54 gnd nmos W='MN10W'   L='MN10L'
MN11  net56   VB4    gnd gnd nmos W='MN11W'   L='MN11L'
MN12  DM_1    VB3    net56 gnd nmos W='MN12W'   L='MN12L'
I0    net1    gnd    'CURRENT_0_BIAS'
C1    net050  VOUT   'CAPACITOR_0'
C2    net050  net2   'CAPACITOR_1'
.ends leung_dfcfc2_pin_3_amp
