* inv_chain

.subckt inv_chain gnd vdd vin vout
MP0  vinb   vin    vdd  vdd  pmos  W='MP0W'  L='MP0L'
MN0  vinb   vin    gnd  gnd  nmos  W='MN0W'  L='MN0L'
MP1  vinbb  vinb   vdd  vdd  pmos  W='MP1W'  L='MP1L'
MN1  vinbb  vinb   gnd  gnd  nmos  W='MN1W'  L='MN1L'
MP2  vinbb  vinb   vdd  vdd  pmos  W='MP2W'  L='MP2L'
MN2  vinbb  vinb   gnd  gnd  nmos  W='MN2W'  L='MN2L'
MP3  vout   vinbb  vdd  vdd  pmos  W='MP3W'  L='MP3L'
MN3  vout   vinbb  gnd  gnd  nmos  W='MN3W'  L='MN3L'
MP4  vout   vinbb  vdd  vdd  pmos  W='MP4W'  L='MP4L'
MN4  vout   vinbb  gnd  gnd  nmos  W='MN4W'  L='MN4L'
MP5  vout   vinbb  vdd  vdd  pmos  W='MP5W'  L='MP5L'
MN5  vout   vinbb  gnd  gnd  nmos  W='MN5W'  L='MN5L'
MP6  vout   vinbb  vdd  vdd  pmos  W='MP6W'  L='MP6L'
MN6  vout   vinbb  gnd  gnd  nmos  W='MN6W'  L='MN6L'
C0   vinb   gnd  'C0'
C1   vinbb  gnd  'C1'
C2   vout   gnd  'C2'
.ends inv_chain