* diode_delay_line

.subckt diode_delay_line gnd vdd vin vout
* first stage
MP0  vin_bar  vin   vdd  vdd  pmos  W='MP0W'  L='MP0L'
MN0  vin_bar  vin   gnd  gnd  nmos  W='MN0W'  L='MN0L'
MN1  vin_bar  VCTRL mn1s gnd  nmos  W='MN1W'  L='MN1L'
MP1  gnd      gnd   mn1s vdd  pmos  W='MP1W'  L='MP1L'
* second stage
MP2  vout  vin_bar  vdd  vdd  pmos  W='MP2W'  L='MP2L'
MN2  vout  vin_bar  gnd  gnd  nmos  W='MN2W'  L='MN2L'
MN3  vout  VCTRL    mn3s gnd  nmos  W='MN3W'  L='MN3L'
MP3  gnd   gnd      mn3s vdd  pmos  W='MP3W'  L='MP3L'
* capacitor
C0   vout  gnd  'C0'
* VCTRL
VCTRL VCTRL 0 'VCTRL'
.ends diode_delay_line