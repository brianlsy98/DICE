* CMOS Inverter with Resistor/Capacitor Load
* DC simulation


* Netlist

.include (MOS_SPEC)

MN0 Vo Vin VSS VSS nmos W=(MN0W) L=(MN0L)

MP0 Vo Vin VDD VDD pmos W=(MP0W) L=(MP0L)

R0  Vo   Vout (R0)
C0  Vout VS   (C0)



* Simulation

.option TEMP=(TEMP)

Vpower  VDD  0  (VDD)
Vgnd    VSS  0  (VSS)
Vinput  Vin  0

.dc Vinput (Vin_min) (Vin_max) (Vin_step)

.control
    run
    wrdata (OUT_PATH) (OUT_DATA)
.endc

.END
