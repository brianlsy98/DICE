* dynamic_latched_comparator

.subckt dynamic_latched_comparator gnd vdd vi_p vi_n vclk vo_p vo_n
MP0  vo_n   vclk    vdd   vdd  pmos  W='MP0W'  L='MP0L'
MP1  vo_n   vo_p    vdd   vdd  pmos  W='MP1W'  L='MP1L'
MP2  vo_p   vo_n    vdd   vdd  pmos  W='MP2W'  L='MP2L'
MP3  vo_p   vclk    vdd   vdd  pmos  W='MP3W'  L='MP3L'
MP4  vg1    vclk    vg2   vdd  pmos  W='MP4W'  L='MP4L'
MN0  va     vin_p   vm    gnd  nmos  W='MN0W'  L='MN0L'
MN1  vo_n   vg1     va    gnd  nmos  W='MN1W'  L='MN1L'
MN2  vb     vin_n   vm    gnd  nmos  W='MN2W'  L='MN2L'
MN3  vo_p   vg2     vb    gnd  nmos  W='MN3W'  L='MN3L'
MN4  vm     vclk    gnd   gnd  nmos  W='MN4W'  L='MN4L'
C0   vo_p   gnd  'C0'
C1   vo_n   gnd  'C1'
C2   vm     gnd  'C2'
.ends dynamic_latched_comparator