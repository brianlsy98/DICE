* NAND

.subckt nand gnd vdd vina vinb vout
MP0  vout  vina  vdd  vdd  pmos  W='MP0W'  L='MP0L'
MP1  vout  vinb  vdd  vdd  pmos  W='MP1W'  L='MP1L'
MN0  mn0d  vina  gnd  gnd  nmos  W='MN0W'  L='MN0L'
MN1  vout  vinb  mn0d  gnd  nmos  W='MN1W'  L='MN1L'
C0   vout  gnd  'C0'
.ends nand