* Simulation for Amplifiers (from AnalogGym)


.include './technology_files/45nm_bulk.txt'
.include './downstream_tasks/opamp_metric_prediction/netlist.cir'


.PARAM supply_voltage = 1.0
.PARAM VCM_ratio = 0.5
.PARAM PARAM_CLOAD = 200.00p 

V1 vdd 0 'supply_voltage'
V2 vss 0 0 

Vindc opin 0 'supply_voltage*VCM_ratio'
Vin signal_in 0 dc 'supply_voltage*VCM_ratio' ac 1 sin('supply_voltage*VCM_ratio' 100m 500)

Lfb opout opout_dc 1T
Cin opout_dc signal_in 1T

* XOP gnda vdda vinn vinp vout
*        |  |     |     |   |
*        |  |     |     |   Output
*        |  |     |     Non-inverting Input
*        |  |      Inverting Input
*        |  Positive Supply
*        Negative Supply 


*    ADM TB   
Xop1 vss vdd opout_dc opin opout  'netlist_name'
Cload1 opout 0 'PARAM_CLOAD'

*    ACM TB    
xop2 vss vdd cm2 cm1 cm3  'netlist_name'
Cload2 cm3 0 'PARAM_CLOAD'
vcmdc cm0 0 'supply_voltage*VCM_ratio'
vcmac1 cm1 cm0 0 ac=1
vcmac2 cm2 cm3 0 ac=1
.meas ac cmrrdc find vdb(cm3) at = 0.1 
.meas ac dcgain find vdb(opout) at = 0.1
.meas ac gain_bandwidth_product when vdb(opout)=0 at = 0.1
.meas ac phase_in_rad find vp(opout) when vdb(opout)=0 at = 0.1

*    PSRR TB
VGNDApsrr gndpsrr 0 0 AC=1
VVDDApsrr vddpsrr 0 'supply_voltage'  AC=1
xop3 vss vddpsrr ppsr1 opin ppsr1  'netlist_name'
Cload3 ppsr1 0 'PARAM_CLOAD'
xop4 gndpsrr vdd npsr1 opin npsr1  'netlist_name'
Cload4 npsr1 0 'PARAM_CLOAD'
.measure ac DCPSRp find vdb(ppsr1) at = 0.1
.measure ac DCPSRn find vdb(npsr1) at = 0.1

*    DC ALL TB
VVDDdc VDDdc 0 'supply_voltage' 
xop5 vss vdddc vout6 opin vout6  'netlist_name'
Cload5 vout6 0 'PARAM_CLOAD'
*    Power meas   
.meas dc Ivdd25 FIND I(VVDDDC) AT=25
.meas dc Power param='-1*Ivdd25*supply_voltage'
*    Vos.meas
.meas dc vout25 FIND V(vout6) AT=25
.meas dc vos25 param = 'vout25-supply_voltage*VCM_ratio'


.control
DC temp  25   26   1
ac dec   10   0.1  1
.endc

.end