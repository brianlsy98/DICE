* AND

.subckt and gnd vdd vina vinb vout
MP0  vout_b  vina    vdd   vdd  pmos  W='MP0W'  L='MP0L'
MP1  vout_b  vinb    vdd   vdd  pmos  W='MP1W'  L='MP1L'
MN0  mn0d    vina    gnd   gnd  nmos  W='MN0W'  L='MN0L'
MN1  vout_b  vinb    mn0d  gnd  nmos  W='MN1W'  L='MN1L'
C0   vout_b  gnd     'C0'
MP2  vout    vout_b  vdd   vdd  pmos  W='MP2W'  L='MP2L'
MN2  vout    vout_b  vdd   vdd  nmos  W='MN2W'  L='MN2L'
C1   vout    gnd     'C1'
.ends and