* Leung_DFCFC2_Pin_3 Amplifier

.subckt leung_dfcfc2_pin_3_amp gnd vdd vinn vinp vout
MP0   vout    net050 vdd vdd pmos W='MP0W'    L='MP0L'
MP1   net049  net1   vdd vdd pmos W='MP1W'    L='MP1L'
MP2   net043  net050 vdd vdd pmos W='MP2W'    L='MP2L'
MP3   net2    net050 vdd vdd pmos W='MP3W'    L='MP3L'
MP4   net050  voutn  vdd vdd pmos W='MP4W'    L='MP4L'
MP5   voutn   voutn  vdd vdd pmos W='MP5W'    L='MP5L'
MP6   net063  vinp   net31 net31 pmos W='MP6W'    L='MP6L'
MP7   dm_2    vinn   net31 net31 pmos W='MP7W'    L='MP7L'
MP8   net31   net1   vdd vdd pmos W='MP8W'    L='MP8L'
MP9   vb3     net1   vdd vdd pmos W='MP9W'    L='MP9L'
MP10  dm_1    net1   vdd vdd pmos W='MP10W'   L='MP10L'
MP11  vb4     net1   vdd vdd pmos W='MP11W'   L='MP11L'
MP12  net1    net1   vdd vdd pmos W='MP12W'   L='MP12L'
MN0   vout    net049 gnd gnd nmos W='MN0W'    L='MN0L'
MN1   net049  net043 gnd gnd nmos W='MN1W'    L='MN1L'
MN2   net043  net043 gnd gnd nmos W='MN2W'    L='MN2L'
MN3   dm_2    vb4    gnd gnd nmos W='MN3W'    L='MN3L'
MN4   voutn   vb3    dm_2 gnd nmos W='MN4W'   L='MN4L'
MN5   net063  vb4    gnd gnd nmos W='MN5W'    L='MN5L'
MN6   net050  vb3    net063 gnd nmos W='MN6W'   L='MN6L'
MN7   net54   vb4    gnd gnd nmos W='MN7W'    L='MN7L'
MN8   net2    vb4    gnd gnd nmos W='MN8W'    L='MN8L'
MN9   vb3     vb3    gnd gnd nmos W='MN9W'    L='MN9L'
MN10  vb4     vb3    net54 gnd nmos W='MN10W'   L='MN10L'
MN11  net56   vb4    gnd gnd nmos W='MN11W'   L='MN11L'
MN12  dm_1    vb3    net56 gnd nmos W='MN12W'   L='MN12L'
I0    net1    gnd    'I0'
C0    net050  vout   'C0'
C1    net050  net2   'C1'
.ends leung_dfcfc2_pin_3_amp
