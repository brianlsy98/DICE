* Yan_AZ_Pin_3 Amplifier

.subckt yan_az_pin_3_amp gnd vdd vinn vinp vout

* PMOS Transistors
MP0   net057  voutn  vdd    vdd    pmos W='MP0W' L='MP0L'
MP1   net078  vb1    vdd    vdd    pmos W='MP1W' L='MP1L'
MP2   vout    net050 vdd    vdd    pmos W='MP2W' L='MP2L'
MP3   net094  net050 vdd    vdd    pmos W='MP3W' L='MP3L'
MP4   net050  voutn  vdd    vdd    pmos W='MP4W' L='MP4L'
MP5   voutn   voutn  vdd    vdd    pmos W='MP5W' L='MP5L'
MP6   net063  vinp   net019 net019 pmos W='MP6W' L='MP6L'
MP7   dm_2    vinn   net019 net019 pmos W='MP7W' L='MP7L'
MP8   net019  vb1    vdd    vdd    pmos W='MP8W' L='MP8L'
MP9   vb4     vb1    vdd    vdd    pmos W='MP9W' L='MP9L'
MP10  vb1     vb1    vdd    vdd    pmos W='MP10W' L='MP10L'

* NMOS Transistors
MN0   net077 dm_2   gnd    gnd nmos W='MN0W' L='MP0L'
MN1   net082 net063 gnd    gnd nmos W='MN1W' L='MN1L'
MN2   vout   net057 gnd    gnd nmos W='MN2W' L='MN2L'
MN3   net094 net051 gnd    gnd nmos W='MN3W' L='MN3L'
MN4   net057 net094 gnd    gnd nmos W='MN4W' L='MN4L'
MN5   dm_2   vb4    gnd    gnd nmos W='MN5W' L='MN5L'
MN6   voutn  net077 dm_2   gnd nmos W='MN6W' L='MN6L'
MN7   net063 vb4    gnd    gnd nmos W='MN7W' L='MN7L'
MN8   net050 net082 net063 gnd nmos W='MN8W' L='MN8L'
MN9   vb4    vb4    gnd    gnd nmos W='MN9W' L='MN9L'

* Current Source
I0 vb1 gnd 'I0'

* Capacitors and Resistors
C1 net051 gnd 'C1'
C0 net063 vout 'C0'
R2 net094 net051 'R2'
R1 net078 net082 'R1'
R0 net078 net077 'R0'

.ends yan_az_pin_3_amp
