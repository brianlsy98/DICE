* Fan_SMC_Pin_3 Amplifier

.subckt fan_smc_pin_3_amp gnd vdd vinn vinp vout
MP0  vout    net050 vdd vdd pmos W='MP0W'   L='MP0L'
MP1  net049  net013 vdd vdd pmos W='MP1W'   L='MP1L'
MP2  net043  net050 vdd vdd pmos W='MP2W'   L='MP2L'
MP3  net050  voutn  vdd vdd pmos W='MP3W'   L='MP3L'
MP4  voutn   voutn  vdd vdd pmos W='MP4W'   L='MP4L'
MP5  net063  vinp   net31 net31 pmos W='MP5W'   L='MP5L'
MP6  dm_2    vinn   net31 net31 pmos W='MP6W'   L='MP6L'
MP7  net31   net013 vdd vdd pmos W='MP7W'   L='MP7L'
MP8  vb3     net013 vdd vdd pmos W='MP8W'   L='MP8L'
MP9  dm_1    net013 vdd vdd pmos W='MP9W'   L='MP9L'
MP10 vb4     net013 vdd vdd pmos W='MP10W'  L='MP10L'
MP11 net013  net013 vdd vdd pmos W='MP11W'  L='MP11L'
MN0  vout    net049 gnd gnd nmos W='MN0W'   L='MN0L'
MN1  net049  net043 gnd gnd nmos W='MN1W'   L='MN1L'
MN2  net043  net043 gnd gnd nmos W='MN2W'   L='MN2L'
MN3  dm_2    vb4    gnd gnd nmos W='MN3W'   L='MN3L'
MN4  voutn   vb3    dm_2 gnd nmos W='MN4W'  L='MN4L'
MN5  net063  vb4    gnd gnd nmos W='MN5W'   L='MN5L'
MN6  net050  vb3    net063 gnd nmos W='MN6W' L='MN6L'
MN7  net54   vb4    gnd gnd nmos W='MN7W'   L='MN7L'
MN8  vb3     vb3    gnd gnd nmos W='MN8W'   L='MN8L'
MN9  vb4     vb3    net54 gnd nmos W='MN9W' L='MN9L'
MN10 net56   vb4    gnd gnd nmos W='MN10W'  L='MN10L'
MN11 dm_1    vb3    net56 gnd nmos W='MN11W' L='MN11L'
I0   net013  gnd    'I0'
C0   net050  vout   'C0'
.ends fan_smc_pin_3_amp
