* capbank_delay_line

.subckt capbank_delay_line gnd vdd vin vout
* inverters
MP0  vin_bar  vin   vdd  vdd  pmos  W='MP0W'  L='MP0L'
MN0  vin_bar  vin   gnd  gnd  nmos  W='MN0W'  L='MN0L'
MP1  vout  vin_bar  vdd  vdd  pmos  W='MP1W'  L='MP1L'
MN1  vout  vin_bar  gnd  gnd  nmos  W='MN1W'  L='MN1L'
* switches
MN2  vin_bar VCTRL0 vc0  gnd  nmos  W='MN2W'  L='MN2L'
MN3  vin_bar VCTRL1 vc1  gnd  nmos  W='MN3W'  L='MN3L'
MN4  vin_bar VCTRL2 vc2  gnd  nmos  W='MN4W'  L='MN4L'
MN5  vin_bar VCTRL3 vc3  gnd  nmos  W='MN5W'  L='MN5L'
MN6  vin_bar VCTRL4 vc4  gnd  nmos  W='MN6W'  L='MN6L'
* capacitors
C0   vc0  gnd  'C0'
C1   vc1  gnd  'C1'
C2   vc2  gnd  'C2'
C3   vc3  gnd  'C3'
C4   vc4  gnd  'C4'
* vctrl
VCTRL0 VCTRL0 0 'VCTRL0'
VCTRL1 VCTRL1 0 'VCTRL1'
VCTRL2 VCTRL2 0 'VCTRL2'
VCTRL3 VCTRL3 0 'VCTRL3'
VCTRL4 VCTRL4 0 'VCTRL4'
.ends capbank_delay_line