* strongarm_latch

.subckt strongarm_latch gnd vdd vi_p vi_n vclk vo_p vo_n
MP0  va    vclk    vdd  vdd  pmos  W='MP0W'  L='MP0L'
MP1  vo_n  vclk    vdd  vdd  pmos  W='MP1W'  L='MP1L'
MP2  vo_n  vo_p    vdd  vdd  pmos  W='MP2W'  L='MP2L'
MP3  vo_p  vo_n    vdd  vdd  pmos  W='MP3W'  L='MP3L'
MP4  vo_p  vclk    vdd  vdd  pmos  W='MP4W'  L='MP4L'
MP5  vb    vclk    vdd  vdd  pmos  W='MP5W'  L='MP5L'
MN0  va    vin_p   vm   gnd  nmos  W='MN0W'  L='MN0L'
MN1  vb    vin_n   vm   gnd  nmos  W='MN1W'  L='MN1L'
MN2  vo_n  vo_p    va   gnd  nmos  W='MN2W'  L='MN2L'
MN3  vo_p  vo_n    vb   gnd  nmos  W='MN3W'  L='MN3L'
MN4  vm    vclk    gnd  gnd  nmos  W='MN4W'  L='MN4L'

C0   vo_p   gnd  'C0'
C1   vo_n   gnd  'C1'
.ends strongarm_latch