* Qu2017_AZC_Pin_3 Amplifier

.subckt qu2017_azc_pin_3_amp gnd vdd vinn vinp vout

* PMOS Transistors
MP0   net057 net055 vdd vdd pmos W='MP0W'  L='MP0L'
MP1   net055 net055 vdd vdd pmos W='MP1W'  L='MP1L'
MP2   net078 vb1     vdd vdd pmos W='MP2W' L='MP2L'
MP3   vout   net050  vdd vdd pmos W='MP3W' L='MP3L'
MP4   net049 vb1     vdd vdd pmos W='MP4W' L='MP4L'
MP5   net094 net050  vdd vdd pmos W='MP5W' L='MP5L'
MP6   net050 voutn   vdd vdd pmos W='MP6W' L='MP6L'
MP7   voutn  voutn   vdd vdd pmos W='MP7W' L='MP7L'
MP8   net063 vinp    net019 net019 pmos W='MP8W'  L='MP8L'
MP9   dm_2   vinn    net019 net019 pmos W='MP9W'  L='MP9L'
MP10  net019 vb1     vdd vdd pmos W='MP10W' L='MP10L'
MP11  vb4    vb1     vdd vdd pmos W='MP11W' L='MP11L'
MP12  vb1    vb1     vdd vdd pmos W='MP12W' L='MP12L'

* NMOS Transistors
MN0   net049 net057 gnd gnd nmos W='MN0W'  L='MN0L'
MN1   net055 net094 gnd gnd nmos W='MN1W'  L='MN1L'
MN2   net077 dm_2   gnd gnd nmos W='MN2W'  L='MN2L'
MN3   net082 net063 gnd gnd nmos W='MN3W'  L='MN3L'
MN4   vout   net049  gnd gnd nmos W='MN4W'  L='MN4L'
MN5   net094 net051 gnd gnd nmos W='MN5W'  L='MN5L'
MN6   net057 net043 gnd gnd nmos W='MN6W'  L='MN6L'
MN7   dm_2   vb4    gnd gnd nmos W='MN7W'  L='MN7L'
MN8   voutn  net077 dm_2 gnd nmos W='MN8W'  L='MN8L'
MN9   net063 vb4    gnd gnd nmos W='MN9W'  L='MN9L'
MN10  net050 net082 net063 gnd nmos W='MN10W' L='MN10L'
MN11  vb4    vb4    gnd gnd nmos W='MN11W' L='MN11L'

* Current Source
I0    vb1    gnd 'I0'

* Capacitors
C2    net043 gnd 'C2'
C1    net051 gnd 'C1'
C0    net063 vout 'C0'

* Resistors
R3    net057 net043 'R3'
R2    net057 net051 'R2'
R1    net078 net082 'R1'
R0    net078 net077 'R0'

.ends qu2017_azc_pin_3_amp
