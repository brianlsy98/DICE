* moscap_delay_line

.subckt moscap_delay_line gnd vdd vin vout
* first stage inv
MP0  vin_bar  vin   vdd  vdd  pmos  W='MP0W'  L='MP0L'
MN0  vin_bar  vin   gnd  gnd  nmos  W='MN0W'  L='MN0L'
* second stage inv
MP1  vout  vin_bar  vdd  vdd  pmos  W='MP1W'  L='MP1L'
MN1  vout  vin_bar  gnd  gnd  nmos  W='MN1W'  L='MN1L'
* switches
MN2  vin_bar  VCTRL0  mn2s  gnd  nmos  W='MN2W'  L='MN2L'
MN3  vin_bar  VCTRL1  mn3s  gnd  nmos  W='MN3W'  L='MN3L'
MN4  vin_bar  VCTRL2  mn4s  gnd  nmos  W='MN4W'  L='MN4L'
* capacitors
MN5  gnd mn2s gnd gnd nmos W='MN5W' L='MN5L'
MN6  gnd mn3s gnd gnd nmos W='MN6W' L='MN6L'
MN7  gnd mn4s gnd gnd nmos W='MN7W' L='MN7L'
C0   vout  gnd  'C0'
* vctrls
VCTRL0 VCTRL0 0 'VCTRL0'
VCTRL1 VCTRL1 0 'VCTRL1'
VCTRL2 VCTRL2 0 'VCTRL2'
.ends moscap_delay_line