* nand_4in

.subckt nand_4in gnd vdd vina vinb vinc vind vout
MP0  vout  vina  vdd   vdd  pmos  W='MP0W'  L='MP0L'
MP1  vout  vinb  vdd   vdd  pmos  W='MP1W'  L='MP1L'
MP2  vout  vinc  vdd   vdd  pmos  W='MP2W'  L='MP2L'
MP3  vout  vind  vdd   vdd  pmos  W='MP3W'  L='MP3L'
MN0  mn0d  vina  gnd   gnd  nmos  W='MN0W'  L='MN0L'
MN1  mn1d  vinb  mn0d  gnd  nmos  W='MN1W'  L='MN1L'
MN2  mn2d  vinc  mn1d  gnd  nmos  W='MN2W'  L='MN2L'
MN3  vout  vind  mn2d  gnd  nmos  W='MN3W'  L='MN3L'
C0   vout  gnd  'C0'
.ends nand_4in