* Yan_AZ_Pin_3 Amplifier

.subckt yan_az_pin_3_amp gnd vdd vinn vinp vout

* PMOS Transistors
MP0   net057 voutn vdd vdd pmos W='MOSFET_0_14_W_BIASCM_PMOS*1' L='MOSFET_0_14_L_BIASCM_PMOS'
MP1   net078 VB1 vdd vdd pmos W='MOSFET_0_14_W_BIASCM_PMOS*1' L='MOSFET_0_14_L_BIASCM_PMOS'
MP2   vout net050 vdd vdd pmos W='MOSFET_13_1_W_gmf2_PMOS*1' L='MOSFET_13_1_L_gmf2_PMOS'
MP3   net094 net050 vdd vdd pmos W='MOSFET_11_1_W_gm2_PMOS*1' L='MOSFET_11_1_L_gm2_PMOS'
MP4   net050 voutn vdd vdd pmos W='MOSFET_0_14_W_BIASCM_PMOS*1' L='MOSFET_0_14_L_BIASCM_PMOS'
MP5   voutn voutn vdd vdd pmos W='MOSFET_0_14_W_BIASCM_PMOS*1' L='MOSFET_0_14_L_BIASCM_PMOS'
MP6   net063 vinp net019 net019 pmos W='MOSFET_9_2_W_gm1_PMOS*1' L='MOSFET_9_2_L_gm1_PMOS'
MP7   DM_2 vinn net019 net019 pmos W='MOSFET_9_2_W_gm1_PMOS*1' L='MOSFET_9_2_L_gm1_PMOS'
MP8   net019 VB1 vdd vdd pmos W='MOSFET_0_14_W_BIASCM_PMOS*1' L='MOSFET_0_14_L_BIASCM_PMOS'
MP9   VB4 VB1 vdd vdd pmos W='MOSFET_0_14_W_BIASCM_PMOS*1' L='MOSFET_0_14_L_BIASCM_PMOS'
MP10  VB1 VB1 vdd vdd pmos W='MOSFET_0_14_W_BIASCM_PMOS*1' L='MOSFET_0_14_L_BIASCM_PMOS'

* NMOS Transistors
MN0   net077 DM_2 gnd gnd nmos W='MOSFET_16_4_W_gm5_NMOS*1' L='MOSFET_16_4_L_gm5_NMOS'
MN1   net082 net063 gnd gnd nmos W='MOSFET_16_4_W_gm5_NMOS*1' L='MOSFET_16_4_L_gm5_NMOS'
MN2   vout net057 gnd gnd nmos W='MOSFET_18_1_W_gm3_NMOS*1' L='MOSFET_18_1_L_gm3_NMOS'
MN3   net094 net051 gnd gnd nmos W='MOSFET_22_1_W_gmb1_NMOS*1' L='MOSFET_22_1_L_gmb1_NMOS'
MN4   net057 net094 gnd gnd nmos W='MOSFET_23_1_W_gmb2_NMOS*1' L='MOSFET_23_1_L_gmb2_NMOS'
MN5   DM_2 VB4 gnd gnd nmos W='MOSFET_19_16_W_BIASCM_NMOS*1' L='MOSFET_19_16_L_BIASCM_NMOS'
MN6   voutn net077 DM_2 gnd nmos W='MOSFET_14_4_W_gm8_NMOS*1' L='MOSFET_14_4_L_gm8_NMOS'
MN7   net063 VB4 gnd gnd nmos W='MOSFET_19_16_W_BIASCM_NMOS*1' L='MOSFET_19_16_L_BIASCM_NMOS'
MN8   net050 net082 net063 gnd nmos W='MOSFET_14_4_W_gm8_NMOS*1' L='MOSFET_14_4_L_gm8_NMOS'
MN9   VB4 VB4 gnd gnd nmos W='MOSFET_19_16_W_BIASCM_NMOS*1' L='MOSFET_19_16_L_BIASCM_NMOS'

* Current Source
I0 VB1 gnd 'CURRENT_1_BIAS'

* Capacitors and Resistors
C1 net051 gnd 'CAPACITOR_0'
C0 net063 vout 'CAPACITOR_1'
R2 net094 net051 'RESISTOR_0'
R1 net078 net082 'RESISTOR_2'
R0 net078 net077 'RESISTOR_1'

.ends yan_az_pin_3_amp
