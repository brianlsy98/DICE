* nor_3in

.subckt nor_3in gnd vdd vina vinb vout
MP0  mp0d  vina  vdd   vdd  pmos  W='MP0W'  L='MP0L'
MP1  mp1d  vinb  mp0d  vdd  pmos  W='MP1W'  L='MP1L'
MP2  vout  vinc  mp1d  vdd  pmos  W='MP2W'  L='MP2L'
MN0  vout  vina  gnd   gnd  nmos  W='MN0W'  L='MN0L'
MN1  vout  vinb  gnd   gnd  nmos  W='MN1W'  L='MN1L'
MN2  vout  vinc  gnd   gnd  nmos  W='MN2W'  L='MN2L'
C0   vout  gnd  'C0'
.ends nor_3in